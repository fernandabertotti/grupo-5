library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sadv1-tb is
end sadv1-tb;

architecture tb of sadv1-tb is
  CONSTANT n_bits : natural := 8;
  signal clk : std_logic := '0';
  
  
