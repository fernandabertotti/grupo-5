--inicializando pasta
